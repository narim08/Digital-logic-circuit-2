module cla4(a, b, ci, s, co); 
  input [3:0] a, b;
  input ci; 
  output [3:0] s; 
  output co;
  wire [3:0] c; 
  
  //full adder module instance
  fa_v2 fa_1(.a(a[0]), .b(b[0]), .ci(ci), .s(s[0]));
  fa_v2 fa_2(.a(a[1]), .b(b[1]), .ci(c[0]), .s(s[1]));
  fa_v2 fa_3(.a(a[2]), .b(b[2]), .ci(c[1]), .s(s[2]));
  fa_v2 fa_4(.a(a[3]), .b(b[3]), .ci(c[2]), .s(s[3]));
  
  //4-bit CLA Block module instance
  clb4 clb4_0(.a(a), .b(b), .ci(ci), .c1(c[0]), .c2(c[1]), .c3(c[2]), .co(co));
  
endmodule
